LIBRARY IEEE; USE IEEE.std_logic_1164.ALL;  USE IEEE.std_logic_unsigned.ALL;  

ENTITY memory1 IS
	GENERIC (blocksize : integer := 4096; segmentsno : integer := 64);
	PORT (
		clk : in std_logic;
		addressbus : IN  STD_LOGIC_VECTOR (11 DOWNTO 0);
		databus : inOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		readmem : in std_logic;
		WriteMem : in std_logic;
		memdataready : OUT std_logic
		);
END memory1;


ARCHITECTURE behavioral OF memory1 IS
	signal data :STD_LOGIC_VECTOR (15 DOWNTO 0); 
	
	--  address 0-127   programs
	--  address 128-134 samples
	--  address 192 -198 data
	
	TYPE mem_TYPE IS ARRAY (0 TO blocksize-1) OF STD_LOGIC_VECTOR (15 DOWNTO 0);   --Data TYPE for a seqment OF memory
	signal mem_array : mem_TYPE:= (
		
		0 =>   "0000011000000000",  -- cwp
		1 =>   "1111110010000000",  -- mil r3 ,128     r3 <= 128;
		2 =>   "0010101100000000",	-- lda r2 , (r3)
		3 =>   "1110100100000000",  -- cmp r2, r1 
		4 =>   "0000100100000100",  -- brc 9
		7 =>   "1111001100000000",  -- jmp 0 
		
		8  =>  "1100100000000000",  -- sub R2-R0-C
		9  =>  "0011111000000000",  -- lda (r3), r2
		10 =>  "0000101000000100",  -- awp 4
		
		
		11 =>  "1111110010000100",  --mil r3 ,132     r3 <= 132;
		12 =>  "0010101100000000",  --lda r2 , (r3)
		13 =>  "1111110011000001",  --mil r3 ,193     r3 <= 193;
		14 =>  "0010011100000000",  --lda r1 , (r3)
		15 =>  "1101011000000000",  --mul r1 , r2
		16 =>  "1011000100000000",  --add r0 , r1
		
		17 =>  "1111110010000101",  --mil r3 ,133     r3 <= 133;
		18 =>  "0010101100000000",  --lda r2 , (r3)
		19 =>  "1111110011000010",  --mil r3 ,194     r3 <= 194;
		20 =>  "0010011100000000",  --lda r1 , (r3)
		21 =>  "1101011000000000",  --mul r1 , r2
		22 =>  "1011000100000000",  --add r0 , r1
		
		23 =>  "1111110010000110",  --mil r3 ,134     r3 <= 134;
		24 =>  "0010101100000000",  --lda r2 , (r3)
		25 =>  "1111110011000011",  --mil r3 ,195     r3 <= 195;
		26 =>  "0010011100000000",  --lda r1 , (r3)
		27 =>  "1101011000000000",  --mul r1 , r2
		28 =>  "1011000100000000",  --add r0 , r1
		
		29 =>  "1111110010000111",  --mil r3 ,135     r3 <= 135;
		30 =>  "0010101100000000",  --lda r2 , (r3)
		31 =>  "1111110011000100",  --mil r3 ,196     r3 <= 196;
		32 =>  "0010011100000000",  --lda r1 , (r3)
		33 =>  "1101011000000000",  --mul r1 , r2
		34 =>  "1011000100000000",  --add r0 , r1
		
		35 =>  "1111110010001000",  --mil r3 ,136     r3 <= 136;
		36 =>  "0010101100000000",  --lda r2 , (r3)
		37 =>  "1111110011000101",  --mil r3 ,197     r3 <= 197;
		38 =>  "0010011100000000",  --lda r1 , (r3)
		39 =>  "1101011000000000",  --mul r1 , r2
		40 =>  "1011000100000000",  --add r0 , r1
		
		41 =>  "1111110010001001",  --mil r3 ,137     r3 <= 137;
		42 =>  "0010011100000000",  --lda r1 , (r3)
		43 =>  "1111110011000110",  --mil r3 ,198     r3 <= 198;
		44 =>  "0010101100000000",  --lda r2 , (r3)
		45 =>  "1101011000000000",  --mul r1 , r2
		46 =>  "1011000100000000",  --add r0 , r1
		
		
		
		47 =>  "1111110010001001",  --mil r3 ,137     r3 <= 137;
		48 =>  "0010011100000000",  --lda r1 , (r3)
		49 =>  "1111110010001010",  --mil r3 ,138     r3 <= 138;
		50 =>  "0011110100000000",  --lda (r3), r1
		
		51 =>  "1111110010001000",  --mil r3 ,136     r3 <= 136;
		52 =>  "0010011100000000",  --lda r1 , (r3)
		53 =>  "1111110010001001",  --mil r3 ,137     r3 <= 137;
		54 =>  "0011110100000000",  --lda (r3), r1
		
		55 =>  "1111110010000111",  --mil r3 ,135     r3 <= 135;
		56 =>  "0010011100000000",  --lda r1 , (r3)
		57 =>  "1111110010001000",  --mil r3 ,136     r3 <= 136;
		58 =>  "0011110100000000",  --lda (r3), r1
		
		59 =>  "1111110010000110",  --mil r3 ,134     r3 <= 134;
		60 =>  "0010011100000000",  --lda r1 , (r3)
		61 =>  "1111110010000111",  --mil r3 ,135     r3 <= 135;
		62 =>  "0011110100000000",  --lda (r3), r1
		
		63 =>  "1111110010000101",  --mil r3 ,133     r3 <= 133;
		64 =>  "0010011100000000",  --lda r1 , (r3)
		65 =>  "1111110010000110",  --mil r3 ,134     r3 <= 134;
		66 =>  "0011110100000000",  --lda (r3), r1
		
		67 =>  "1111110010000100",  --mil r3 ,132     r3 <= 132;
		68 =>  "0010011100000000",  --lda r1 , (r3)
		69 =>  "1111110010000101",  --mil r3 ,133     r3 <= 133;
		70 =>  "0011110100000000",  --lda (r3), r1
		
		71 =>  "1111110010000011",  --mil r3 ,131     r3 <= 131;
		72 =>  "0010011100000000",  --lda r1 , (r3)
		73 =>  "1111110010000100",  --mil r3 ,132     r3 <= 132;
		74 =>  "0011110100000000",  --lda (r3), r1
		
		75 =>  "1111110010000010",  --mil r3 ,130     r3 <= 130;
		76 =>  "0010011100000000",  --lda r1 , (r3)
		77 =>  "1111110010000011",  --mil r3 ,131     r3 <= 131;
		78 =>  "0011110100000000",  --lda (r3), r1
		
		79 =>  "1111110010000001",  --mil r3 ,129     r3 <= 129;
		80 =>  "0010011100000000",  --lda r1 , (r3)
		81 =>  "1111100000000000",  --mil r2 ,0       r2 <= 0;
		82 =>  "0011111000000000",  --lda (r3), r2
		83 =>  "1111110010000010",  --mil r3 ,130     r3 <= 130;
		84 =>  "0011110100000000",  --lda (r3), r1
		85 =>  "1111110010100000",  --mil r3 ,160     r3 <= 160;
		86 =>  "0011110000000000",  --lda (r3), r0
		87 =>  "1111000000000000",  --mil r0 ,0       r2 <= 0;
		88 =>  "1111000100000000",  --miH r0 ,0       r2 <= 0;
		
		
		89 =>  "0000101000001000",  -- awp 8
		90 =>  "1111110010100000",  --mil r3 ,160   r3 <= 160;
		91 =>  "0010011100000000",  --lda r1 , (r3)
		92 =>  "1111100100010000",  --mih r2 ,16    r3 <= 4096;
		93 =>  "0011100100000000",  --lda (r2), r1
		94 =>  "0000010000000000",  --szf   carry <= '1';
		95 =>  "1011100000000000",  --add r2 , r0
		96 =>  "0000101000001000",  -- awp 8
		97 =>  "1111111100000000",  -- jpa r3, 0
		
		
		-- address 128-134 samples
		128 => "0000000000000100",
		129 => "0000000000011101",
		130 => "0000000000001011",
		131 => "0000000000010101",
		132 => "0000000000001001",
		
		
		--  address 192 -198 data
		--192 => "0000000000000110",
		193 => "0000000000010111",
		194 => "0000000000011101",
		195 => "0000000000010110",
		196 => "0000000000011001",
		197 => "0000000000011010",
		198 => "0000000000010101",
		
		
	others => (others => '0'));
	
	
BEGIN
	memdataready <= '1';
	databus <= data when readmem='1' else (others => 'Z');
	
	process	(clk)
	begin
		if (WriteMem='1') and (clk='1' and clk'event) then
			mem_array (conv_integer (addressbus)) <=  databus;
		end if;
	end process;
	
	
	process	(addressbus, ReadMem)
	begin
		if (ReadMem='1') then
			data <= mem_array (conv_integer (addressbus));
		end if;
	end process;
	
END behavioral;
