LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY REGISTERFILE IS
	PORT (
		INPUT : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		CLK, RST : IN STD_LOGIC;
		BASE : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		LADDR, RADDR : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		RFLWRITE, RFHWRITE : IN STD_LOGIC;
		LOUT, ROUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
		);
END REGISTERFILE;

ARCHITECTURE DATAFLOW OF REGISTERFILE IS 
	
	SIGNAL LADDRESS, RADDRESS : STD_LOGIC_VECTOR (5 DOWNTO 0);
	TYPE MEMTYPE IS ARRAY (0 TO 23) OF STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL MEMORYFILE : MEMTYPE;
	
BEGIN
	LADDRESS <= BASE + LADDR;
	RADDRESS <= BASE + RADDR;
	
	LOUT <= MEMORYFILE (CONV_INTEGER(LADDRESS));
	ROUT <= MEMORYFILE (CONV_INTEGER(RADDRESS));
	
	PROCESS (CLK, RST)
	BEGIN 
		IF RST='1' THEN
			MEMORYFILE <= (OTHERS => (OTHERS => '0'));
		ELSIF (CLK = '1') THEN
			IF (RFLWRITE = '1') THEN
				MEMORYFILE (CONV_INTEGER (LADDRESS)) (7 DOWNTO 0) <= INPUT (7 DOWNTO 0);
			END IF;
			IF (RFHWRITE = '1') THEN
				MEMORYFILE (CONV_INTEGER (LADDRESS)) (15 DOWNTO 8) <= INPUT (15 DOWNTO 8);
			END IF;
		END IF;
	END PROCESS;
	
END DATAFLOW;