LIBRARY IEEE;
 USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PROGRAMCOUNTER IS
	PORT (
		ENABLEPC : IN STD_LOGIC;
		INPUT : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		CLK : IN STD_LOGIC;
		OUTPUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
		);
END PROGRAMCOUNTER;

ARCHITECTURE DATAFLOW OF PROGRAMCOUNTER IS
BEGIN
	
	PROCESS (CLK)
	BEGIN
		IF (CLK = '1') THEN
			IF (ENABLEPC = '1') THEN
				OUTPUT <= INPUT;
			END IF;
		END IF;
	END PROCESS;
	
END DATAFLOW;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ADDRESSLOGIC IS
	PORT (
		PCSIDE, RSIDE : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		ISIDE : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		ALOUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		RESETPC, PCPLUSI, PCPLUS1, RPLUSI, RPLUS0 : IN STD_LOGIC
		);
END ADDRESSLOGIC;

ARCHITECTURE DATAFLOW OF ADDRESSLOGIC IS
	CONSTANT ONE   : STD_LOGIC_VECTOR (4 DOWNTO 0) := "10000";
	CONSTANT TWO   : STD_LOGIC_VECTOR (4 DOWNTO 0) := "01000";
	CONSTANT THREE : STD_LOGIC_VECTOR (4 DOWNTO 0) := "00100";
	CONSTANT FOUR  : STD_LOGIC_VECTOR (4 DOWNTO 0) := "00010";
	CONSTANT FIVE  : STD_LOGIC_VECTOR (4 DOWNTO 0) := "00001";
	
BEGIN
	
	PROCESS (PCSIDE, RSIDE, ISIDE, RESETPC, PCPLUSI, PCPLUS1, RPLUSI, RPLUS0)
		VARIABLE TEMP : STD_LOGIC_VECTOR (4 DOWNTO 0);
	BEGIN
		TEMP := (RESETPC & PCPLUSI & PCPLUS1 & RPLUSI & RPLUS0 );
		CASE TEMP IS
			WHEN ONE  => ALOUT <= (OTHERS=>'0');
			WHEN TWO  => ALOUT <= PCSIDE + ISIDE;
			WHEN THREE => ALOUT <= PCSIDE + 1;
			WHEN FOUR  => ALOUT <= RSIDE + ISIDE;
			WHEN FIVE  => ALOUT <= RSIDE;
			WHEN OTHERS => ALOUT <= PCSIDE;
		END CASE;
	END PROCESS;
	
END DATAFLOW;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ADDRESSINGUNIT IS
	PORT (
		RSIDE : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		ISIDE : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		ADDRESS : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		CLK, RESETPC, PCPLUSI, PCPLUS1, RPLUSI, RPLUS0, ENABLEPC : IN STD_LOGIC
		);
END ADDRESSINGUNIT;

ARCHITECTURE DATAFLOW OF ADDRESSINGUNIT IS
	COMPONENT PC
		PORT (
			ENABLEPC : IN STD_LOGIC;
			INPUT : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			CLK : IN STD_LOGIC;
			OUTPUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
			);
	END COMPONENT;
	FOR ALL : PC USE ENTITY WORK.PROGRAMCOUNTER (DATAFLOW);
	
	COMPONENT AL
		PORT (
			PCSIDE, RSIDE : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			ISIDE : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			ALOUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			RESETPC, PCPLUSI, PCPLUS1, RPLUSI, RPLUS0 : IN STD_LOGIC
			);
	END COMPONENT;
	FOR ALL : AL USE ENTITY WORK.ADDRESSLOGIC (DATAFLOW);
	
	SIGNAL PCOUT : STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL ADDRESSSIGNAL : STD_LOGIC_VECTOR (15 DOWNTO 0);
	
BEGIN
	ADDRESS <= ADDRESSSIGNAL;
	
	L1 : PC PORT MAP (ENABLEPC, ADDRESSSIGNAL, CLK, PCOUT);
	L2 : AL PORT MAP (PCOUT, RSIDE, ISIDE, ADDRESSSIGNAL, RESETPC, PCPLUSI, PCPLUS1, RPLUSI, RPLUS0);
END DATAFLOW;
