------- Saye Data Pqath
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DATAPATH IS
	PORT (
		CLK : IN STD_LOGIC;
		DATABUS : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		ADDRESSBUS : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		RESETPC, PCPLUSI, PCPLUS1, RPLUSI, RPLUS0, RS_ON_ADDRESSUNITRSIDE, RD_ON_ADDRESSUNITRSIDE, ENABLEPC, 
		B15TO0, 
		AADDB, ASUBB, AMULB, ACMPB, RFLWRITE, RFHWRITE, WPRESET,
		WPADD, IRLOAD, SRLOAD, ADDRESS_ON_DATABUS, ALU_ON_DATABUS, IR_ON_LOPNDBUS, IR_ON_HOPNDBUS, 
		RFRIGHT_ON_OPNDBUS, CSET, CRESET, ZSET, ZRESET, SHADOW : IN STD_LOGIC;
		INSTRUCTION : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		COUT, ZOUT, SHADOWEN : OUT STD_LOGIC
		);
END DATAPATH;

ARCHITECTURE DATAFLOW OF DATAPATH IS
	COMPONENT AU
		PORT (
			RSIDE : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			ISIDE : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			ADDRESS : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			CLK, RESETPC, PCPLUSI, PCPLUS1, RPLUSI, RPLUS0, ENABLEPC : IN STD_LOGIC
			);
	END COMPONENT;
	FOR ALL : AU USE ENTITY WORK.ADDRESSINGUNIT (DATAFLOW);
	
	COMPONENT ALU
		PORT (
			A, B : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			B15TO0,
			--AANDB, AORB, NOTB, SHLB, SHRB,
			AADDB, ASUBB, AMULB, ACMPB : IN STD_LOGIC;
			ALUOUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			CIN : IN STD_LOGIC;
			ZOUT, COUT : OUT STD_LOGIC
			);
	END COMPONENT;
	FOR ALL : ALU USE ENTITY WORK.ARITHMETICUNIT (DATAFLOW);
	
	COMPONENT RF
		PORT (
			INPUT : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			CLK,RST : IN STD_LOGIC;
			BASE : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
			LADDR, RADDR : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			RFLWRITE, RFHWRITE : IN STD_LOGIC;
			LOUT, ROUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
			);
	END COMPONENT;
	FOR ALL : RF USE ENTITY WORK.REGISTERFILE (DATAFLOW);
	
	COMPONENT IR
		PORT (
			INPUT : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			IRLOAD, CLK : IN STD_LOGIC;
			OUTPUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
			);
	END COMPONENT;
	FOR ALL : IR USE ENTITY WORK.INSTRUNCTIONREGISTER (DATAFLOW);
	
	COMPONENT SR
		PORT (
			CIN, ZIN, SRLOAD, CLK, CSET, CRESET, ZSET, ZRESET : IN STD_LOGIC;
			COUT, ZOUT : OUT STD_LOGIC
			);
	END COMPONENT;
	FOR ALL : SR USE ENTITY WORK.STATUSREGISTER (DATAFLOW);
	
	COMPONENT WP
		PORT (
			INPUT : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
			CLK, WPRESET, WPADD : IN STD_LOGIC;
			OUTPUT : OUT STD_LOGIC_VECTOR (5 DOWNTO 0)
			);
	END COMPONENT;
	FOR ALL : WP USE ENTITY WORK.WINDOWPOINTER (DATAFLOW);
	
	SIGNAL RIGHT, LEFT, OPNDBUS, ALUOUT, IROUT, ADDRESS, ADDRESSUNITRSIDEBUS : STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL SRCIN, SRZIN, SRZOUT, SRCOUT : STD_LOGIC; 
	SIGNAL WPOUT : STD_LOGIC_VECTOR (5 DOWNTO 0);
	SIGNAL LADDR, RADDR : STD_LOGIC_VECTOR (1 DOWNTO 0);
	
BEGIN
	
	ADDRESSINGUNIT : AU PORT MAP (
		ADDRESSUNITRSIDEBUS, IROUT (7 DOWNTO 0), ADDRESS, CLK, RESETPC, PCPLUSI, PCPLUS1, RPLUSI, RPLUS0, ENABLEPC
		);
	
	ARITHMETICUNIT : ALU PORT MAP (
		LEFT, OPNDBUS, B15TO0,
		--AANDB, AORB, NOTB, SHLB, SHRB, 
		AADDB, ASUBB, AMULB, ACMPB, 
		ALUOUT, SRCOUT, SRZIN, SRCIN
		);
	
	REGISTERFILE : RF PORT MAP (
		DATABUS, CLK, RESETPC, WPOUT, LADDR, RADDR, RFLWRITE, RFHWRITE, LEFT, RIGHT
		);
	
	INSTRUNCTIONREGISTER : IR PORT MAP (DATABUS, IRLOAD, CLK, IROUT);
	
	STATUSREGISTER : SR PORT MAP (SRCIN, SRZIN, SRLOAD, CLK, CSET, CRESET, ZSET, ZRESET, SRCOUT, SRZOUT);
	
	WINDOWPOINTER : WP PORT MAP (IROUT (5 DOWNTO 0), CLK, WPRESET, WPADD, WPOUT);
	
	ADDRESSUNITRSIDEBUS <= 
	RIGHT WHEN RS_ON_ADDRESSUNITRSIDE='1' ELSE LEFT WHEN RD_ON_ADDRESSUNITRSIDE='1' ELSE (OTHERS=>'Z');
	
	ADDRESSBUS <= ADDRESS;
	
	DATABUS <= ADDRESS WHEN ADDRESS_ON_DATABUS = '1' ELSE ALUOUT WHEN ALU_ON_DATABUS = '1' ELSE (OTHERS=>'Z');
	
	OPNDBUS (7 DOWNTO 0) <= IROUT (7 DOWNTO 0) WHEN IR_ON_LOPNDBUS = '1' ELSE (OTHERS=>'Z');
	
	OPNDBUS (15 DOWNTO 8) <= IROUT (7 DOWNTO 0) WHEN IR_ON_HOPNDBUS = '1' ELSE (OTHERS=>'Z');
	
	OPNDBUS <= RIGHT WHEN RFRIGHT_ON_OPNDBUS = '1' ELSE (OTHERS=>'Z');
	
	ZOUT <= SRZOUT;
	
	COUT <= SRCOUT;
	
	INSTRUCTION <= IROUT(15 DOWNTO 8) WHEN SHADOW='0' ELSE IROUT(7 DOWNTO 0);
	
	SHADOWEN <= '0' WHEN IROUT (7 DOWNTO 0)="00001111" ELSE '1';
	
	LADDR <= IROUT (11 DOWNTO 10) WHEN SHADOW='0' ELSE IROUT (3 DOWNTO 2);
	
	RADDR <= IROUT (9 DOWNTO 8) WHEN SHADOW='0' ELSE IROUT (1 DOWNTO 0);
	
END DATAFLOW;
