
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY STATUSREGISTER IS
	PORT (
		CIN, ZIN, SRLOAD, CLK, CSET, CRESET, ZSET, ZRESET : IN STD_LOGIC;
		COUT, ZOUT : OUT STD_LOGIC
		);
END STATUSREGISTER;

ARCHITECTURE DATAFLOW OF STATUSREGISTER IS
BEGIN
	
	PROCESS (CLK)
	BEGIN
		IF (CLK = '1') THEN
			IF (SRLOAD = '1') THEN
				COUT <= CIN;
				ZOUT <= ZIN;
			ELSIF (CSET='1') THEN
				COUT <= '1';
			ELSIF (CRESET='1') THEN
				COUT <= '0';
			ELSIF (ZSET='1') THEN
				ZOUT <= '1';
			ELSIF (ZRESET='1') THEN
				ZOUT <= '0';
			END IF;
		END IF;
	END PROCESS;
	
END DATAFLOW;