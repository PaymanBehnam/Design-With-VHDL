							  
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 

ENTITY M1X1 IS
	PORT (XI, YI, PI, CI : IN STD_LOGIC; 
		XO, YO, PO, CO : OUT STD_LOGIC);
END M1X1;
ARCHITECTURE BITWISE OF M1X1 IS
	SIGNAL XY : STD_LOGIC;
BEGIN	   
	XY <= XI AND YI;
	CO <= (PI AND XY) OR (PI AND CI) OR (XY AND CI);
	PO <= PI XOR XY XOR CI;
	XO <= XI;
	YO <= YI;
END BITWISE;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 

ENTITY MULT_8BY8 IS
	PORT (X, Y : IN STD_LOGIC_VECTOR (7 DOWNTO 0); 
		Z : OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END MULT_8BY8;   

ARCHITECTURE BITWISE OF MULT_8BY8 IS 
	
	COMPONENT M1X1 
		PORT (XI, YI, PI, CI : IN STD_LOGIC; 
			XO, YO, PO, CO : OUT STD_LOGIC); 
	END COMPONENT; 
	
	TYPE PAIR IS ARRAY (8 DOWNTO 0, 8 DOWNTO 0) OF STD_LOGIC;
	SIGNAL XV, YV, CV, PV : PAIR;
	
BEGIN 
	
	ROWS : FOR I IN X'RANGE GENERATE
		COLS : FOR J IN Y'RANGE GENERATE
			CELL : M1X1 PORT MAP (XV (I, J), YV (I, J), PV (I, J+1), CV (I, J), XV (I, J+1), YV (I+1, J), PV (I+1, J), CV (I, J+1));
		END GENERATE;
	END GENERATE; 
	
	SIDES : FOR I IN X'RANGE GENERATE
		XV (I, 0) <= X (I);
		CV (I, 0) <= '0';
		PV (0, I+1) <= '0';
		PV (I+1, X'LENGTH) <= CV (I, X'LENGTH);
		YV (0, I) <= Y (I);
		Z (I) <= PV (I+1, 0);
		Z (I+X'LENGTH) <= PV (X'LENGTH, I+1);
	END GENERATE;    
	
END BITWISE;