----------------------------
--SAYEH TESTBENCH
----------------------------
LIBRARY IEEE; USE IEEE.STD_LOGIC_1164.ALL; USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TESTSAYEH IS  END TESTSAYEH;

ARCHITECTURE DATAFLOW OF TESTSAYEH IS
	SIGNAL CLK : STD_LOGIC := '0';
	SIGNAL READIO, WRITEIO, EXTERNALRESET, MEMDATAREADY : STD_LOGIC;
	SIGNAL READMEM, WRITEMEM, READMEM_IN, WRITEMEM_IN, READMEM_OUT, WRITEMEM_OUT : STD_LOGIC;
	SIGNAL ADDRESSBUS_CPU, ADDRESSBUS_fir_in, ADDRESSBUS_MEMORY, DATABUS : STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL ADDRESSBUS_MEM : STD_LOGIC_VECTOR (11 DOWNTO 0);
	SIGNAL ADDR_INT : INTEGER;
	
	
	SIGNAL REQUEST1, REQUEST2 : STD_LOGIC;
	SIGNAL READ_OUT, WR_OUT : STD_LOGIC;
	signal MEMREADY_OUT1, MEMREADY_OUT2 : std_logic;
	signal wr_mem_FIR_IN, REQUEST_FIR_IN : std_logic;
BEGIN
	
	CLK <= NOT (CLK) AFTER 5 NS WHEN NOW<1000000 NS ELSE CLK;
	EXTERNALRESET <= '1', '0' AFTER 7 NS;
	
	PROCESSOR : ENTITY WORK.SAYEH(DATAFLOW)  PORT MAP  (
		CLK => CLK,
		READMEM => READMEM,
		WRITEMEM => WRITEMEM,
		READIO => READIO,
		WRITEIO => WRITEIO,
		DATABUS => DATABUS,
		ADDRESSBUS => ADDRESSBUS_CPU,
		EXTERNALRESET => EXTERNALRESET,
		MEMDATAREADY => MEMREADY_OUT1
		);
	
	MEMORY_IN : ENTITY WORK.MEMORY1 (BEHAVIORAL)
	PORT MAP (
		CLK => CLK,
		ADDRESSBUS => ADDRESSBUS_MEM,
		DATABUS => DATABUS,
		READMEM => READMEM_IN,
		WRITEMEM => WRITEMEM_IN,
		MEMDATAREADY => MEMDATAREADY
		);
	
	MEMORY_OUT : ENTITY WORK.MEMORY2 (BEHAVIORAL)
	PORT MAP (
		CLK => CLK,
		ADDRESSBUS => ADDRESSBUS_MEM,
		DATABUS => DATABUS,
		READMEM => READMEM_OUT,
		WRITEMEM => WRITEMEM_OUT,
		MEMDATAREADY => MEMDATAREADY
		);
	
	DMA_MODEL :ENTITY WORK.DMA (DATAFLOW)
	PORT MAP (
		RST => EXTERNALRESET,
		CLK => CLK,
		ADDR_IN1 => ADDRESSBUS_CPU,
		ADDR_IN2 => ADDRESSBUS_fir_in,
		ADDR_OUT => ADDRESSBUS_MEMORY,
		READ_IN1 => READMEM,
		READ_IN2 => '0',
		READ_OUT => READ_OUT,
		WR_IN1 => WRITEMEM,
		WR_IN2 => wr_mem_FIR_IN,
		WR_OUT => WR_OUT,
		REQUEST1 => REQUEST1,
		REQUEST2 => REQUEST_FIR_IN,
		MEMREADY_IN => '1',
		MEMREADY_OUT1 => MEMREADY_OUT1,
		MEMREADY_OUT2 => MEMREADY_OUT2
		);
	
	FIR_IN :entity work.fir_input(behav)
	port map (
		RST => EXTERNALRESET,
		CLK => CLK,
		ADDR_OUT => ADDRESSBUS_fir_in,
		DATAOUT => DATABUS,
		SEND => MEMREADY_OUT2,
		WR => wr_mem_FIR_IN,
		REQUEST => REQUEST_FIR_IN
		);
	
	REQUEST1 <= READMEM OR WRITEMEM;
	
	ADDRESSBUS_MEM <= ADDRESSBUS_MEMORY (11 DOWNTO 0) AFTER 1 NS;
	ADDR_INT <= CONV_INTEGER (ADDRESSBUS_MEMORY);
	READMEM_IN  <= READ_OUT  WHEN (ADDR_INT < 4096 ) ELSE '0';
	WRITEMEM_IN <= WR_OUT WHEN (ADDR_INT < 4096 ) ELSE '0';
	
	READMEM_OUT  <= READ_OUT  WHEN (ADDR_INT > 4095 ) ELSE '0';
	WRITEMEM_OUT <= WR_OUT WHEN (ADDR_INT > 4095 ) ELSE '0';
	
END DATAFLOW;