-- Saye Processor

LIBRARY IEEE; USE IEEE.STD_LOGIC_1164.ALL; USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SAYEH IS
	PORT (
		CLK : IN STD_LOGIC;
		READMEM, WRITEMEM, READIO, WRITEIO : OUT STD_LOGIC;
		DATABUS : INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		ADDRESSBUS : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		EXTERNALRESET, MEMDATAREADY : IN STD_LOGIC
		);
END SAYEH;

ARCHITECTURE DATAFLOW OF SAYEH IS
	
	SIGNAL INSTRUCTION : STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL RESETPC, PCPLUSI, PCPLUS1, RPLUSI, RPLUS0, RS_ON_ADDRESSUNITRSIDE, RD_ON_ADDRESSUNITRSIDE,
		ENABLEPC, B15TO0, BLEAST, AADDB, ASUBB, AMULB, ACMPB, 
		RFLWRITE, RFHWRITE, RFZEROLEFT, RFZERORIGHT, WPRESET, WPADD, IRLOAD, SRLOAD,
		ADDRESS_ON_DATABUS, ALU_ON_DATABUS, IR_ON_LOPNDBUS, IR_ON_HOPNDBUS, RFRIGHT_ON_OPNDBUS,
	CSET, CRESET, ZSET, ZRESET, SHADOW, CFLAG, ZFLAG, SHADOWEN : STD_LOGIC; 
	
BEGIN
	
	DP :ENTITY WORK.DATAPATH
	PORT MAP (
		CLK => CLK,
		DATABUS => DATABUS,
		ADDRESSBUS => ADDRESSBUS,
		RESETPC => RESETPC,
		PCPLUSI => PCPLUSI,
		PCPLUS1 => PCPLUS1,
		RPLUSI => RPLUSI,
		RPLUS0 => RPLUS0,
		RS_ON_ADDRESSUNITRSIDE => RS_ON_ADDRESSUNITRSIDE,
		RD_ON_ADDRESSUNITRSIDE => RD_ON_ADDRESSUNITRSIDE,
		ENABLEPC => ENABLEPC,
		B15TO0 => B15TO0,
		AADDB => AADDB,
		ASUBB => ASUBB,
		AMULB => AMULB,
		ACMPB => ACMPB,
		RFLWRITE => RFLWRITE,
		RFHWRITE => RFHWRITE,
		WPRESET => WPRESET,
		WPADD => WPADD,
		IRLOAD => IRLOAD,
		SRLOAD => SRLOAD,
		ADDRESS_ON_DATABUS => ADDRESS_ON_DATABUS,
		ALU_ON_DATABUS => ALU_ON_DATABUS,
		IR_ON_LOPNDBUS => IR_ON_LOPNDBUS,
		IR_ON_HOPNDBUS => IR_ON_HOPNDBUS,
		RFRIGHT_ON_OPNDBUS => RFRIGHT_ON_OPNDBUS,
		CSET => CSET,
		CRESET => CRESET,
		ZSET => ZSET,
		ZRESET => ZRESET,
		SHADOW => SHADOW,
		INSTRUCTION => INSTRUCTION,
		COUT => CFLAG,
		ZOUT => ZFLAG,
		SHADOWEN => SHADOWEN
		);
	
	CONTROLLER : ENTITY WORK.CONTROLLER	
	PORT MAP (
		EXTERNALRESET => EXTERNALRESET,
		CLK => CLK,
		RESETPC => RESETPC,
		PCPLUSI => PCPLUSI,
		PCPLUS1 => PCPLUS1,
		RPLUSI => RPLUSI,
		RPLUS0 => RPLUS0,
		RS_ON_ADDRESSUNITRSIDE => RS_ON_ADDRESSUNITRSIDE,
		RD_ON_ADDRESSUNITRSIDE => RD_ON_ADDRESSUNITRSIDE,
		ENABLEPC => ENABLEPC,
		B15TO0 => B15TO0,
		AADDB => AADDB,
		ASUBB => ASUBB,
		AMULB => AMULB,
		ACMPB => ACMPB,
		RFLWRITE => RFLWRITE,
		RFHWRITE => RFHWRITE,
		WPRESET => WPRESET,
		WPADD => WPADD,
		IRLOAD => IRLOAD,
		SRLOAD => SRLOAD,
		ADDRESS_ON_DATABUS => ADDRESS_ON_DATABUS,
		ALU_ON_DATABUS => ALU_ON_DATABUS,
		IR_ON_LOPNDBUS => IR_ON_LOPNDBUS,
		IR_ON_HOPNDBUS => IR_ON_HOPNDBUS,
		RFRIGHT_ON_OPNDBUS => RFRIGHT_ON_OPNDBUS,
		READMEM => READMEM,
		WRITEMEM => WRITEMEM,
		CSET => CSET,
		CRESET => CRESET,
		ZSET => ZSET,
		ZRESET => ZRESET,
		SHADOW => SHADOW,
		INSTRUCTION => INSTRUCTION,
		CFLAG => CFLAG,
		ZFLAG => ZFLAG,
		MEMDATAREADY => MEMDATAREADY,
		SHADOWEN => SHADOWEN
		);
	
END DATAFLOW;


