
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ARITHMETICUNIT IS
	PORT (
		A, B : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		B15TO0, 
		--AANDB, AORB, NOTB, SHLB, SHRB,
		AADDB, ASUBB, AMULB, ACMPB : IN STD_LOGIC;
		ALUOUT : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		CIN : IN STD_LOGIC;
		ZOUT, COUT : OUT STD_LOGIC
		);
END ARITHMETICUNIT;

ARCHITECTURE DATAFLOW OF ARITHMETICUNIT IS
	COMPONENT MULT 
		PORT (
			X, Y : IN STD_LOGIC_VECTOR (7 DOWNTO 0); 
			Z : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
			);
	END COMPONENT;
	FOR ALL : MULT USE ENTITY WORK.MULT_8BY8 (BITWISE);
	
	CONSTANT B15TO0H : STD_LOGIC_VECTOR (9 DOWNTO 0) := "1000000000";
	CONSTANT AANDBH  : STD_LOGIC_VECTOR (9 DOWNTO 0) := "0100000000";
	CONSTANT AORBH   : STD_LOGIC_VECTOR (9 DOWNTO 0) := "0010000000";
	CONSTANT NOTBH   : STD_LOGIC_VECTOR (9 DOWNTO 0) := "0001000000";
	CONSTANT SHLBH   : STD_LOGIC_VECTOR (9 DOWNTO 0) := "0000100000";
	CONSTANT SHRBH   : STD_LOGIC_VECTOR (9 DOWNTO 0) := "0000010000";
	CONSTANT AADDBH  : STD_LOGIC_VECTOR (9 DOWNTO 0) := "0000001000";
	CONSTANT ASUBBH  : STD_LOGIC_VECTOR (9 DOWNTO 0) := "0000000100";
	CONSTANT AMULBH  : STD_LOGIC_VECTOR (9 DOWNTO 0) := "0000000010";
	CONSTANT ACMPBH  : STD_LOGIC_VECTOR (9 DOWNTO 0) := "0000000001";
	SIGNAL ALUOUTSIGNAL, PRODUCT : STD_LOGIC_VECTOR (15 DOWNTO 0);
	
BEGIN
	--PROCESS (A, B, B15TO0, AANDB, AORB, NOTB, SHLB, SHRB, AADDB, ASUBB, AMULB, CIN, ALUOUTSIGNAL, PRODUCT, ACMPB)--SIGNAL, PRODUCT ARE ADDED
	PROCESS (A, B, B15TO0, AADDB, ASUBB, AMULB, CIN, ALUOUTSIGNAL, PRODUCT, ACMPB)--SIGNAL, PRODUCT ARE ADDED
		VARIABLE TEMP :  STD_LOGIC_VECTOR (9 DOWNTO 0);
		VARIABLE SUM :  STD_LOGIC_VECTOR (16 DOWNTO 0);
		VARIABLE SUB :  STD_LOGIC_VECTOR (16 DOWNTO 0);
	BEGIN
		ZOUT <= '0';
		COUT <= '0';
		ALUOUTSIGNAL <= (OTHERS=>'0');
		--TEMP := (B15TO0, AANDB, AORB, NOTB, SHLB, SHRB, AADDB, ASUBB, AMULB, ACMPB);
		TEMP := (B15TO0, '0', '0', '0', '0', '0', AADDB, ASUBB, AMULB, ACMPB);
		SUM := ("0"&A) + B + CIN ;
		SUB := ("0"&A) - B - CIN;
		
		CASE TEMP IS
			WHEN B15TO0H => ALUOUTSIGNAL <= B;
			WHEN AADDBH  => ALUOUTSIGNAL <= SUM (15 DOWNTO 0);COUT <= SUM (16);
			WHEN ASUBBH  => ALUOUTSIGNAL <= SUB (15 DOWNTO 0);COUT <= SUB (16);
			WHEN AMULBH  => ALUOUTSIGNAL <= PRODUCT; --A (7 DOWNTO 0) * B (7 DOWNTO 0);
			WHEN ACMPBH  => ALUOUTSIGNAL <= (OTHERS=>'1');
			IF (A>B) THEN
				COUT <= '1';
			ELSE
				COUT <= '0';
			END IF;
			
			IF (A=B) THEN
				ZOUT <= '1';
			ELSE
				ZOUT <= '0';
			END IF;
			WHEN OTHERS => ALUOUTSIGNAL <= (OTHERS=>'0');
		END CASE;
		
		IF (ALUOUTSIGNAL = "0000000000000000") THEN
			ZOUT <= '1';
		END IF;
		
	END PROCESS;
	
	L1 : MULT PORT MAP (A (7 DOWNTO 0), B (7 DOWNTO 0), PRODUCT);
	
	ALUOUT <= ALUOUTSIGNAL;
	
END DATAFLOW;
