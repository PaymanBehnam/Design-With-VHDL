LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY WINDOWPOINTER IS
	PORT (
		INPUT : IN STD_LOGIC_VECTOR (5 DOWNTO 0);
		CLK, WPRESET, WPADD : IN STD_LOGIC;
		OUTPUT : OUT STD_LOGIC_VECTOR (5 DOWNTO 0)
		);
END WINDOWPOINTER;

ARCHITECTURE DATAFLOW OF WINDOWPOINTER IS
	SIGNAL OUTPUTSIGNAL : STD_LOGIC_VECTOR (5 DOWNTO 0);
	
BEGIN
	
	PROCESS (CLK)
	BEGIN
		IF (CLK = '1') THEN
			IF (WPRESET = '1') THEN
				OUTPUTSIGNAL <= (OTHERS => '0');
			ELSIF (WPADD = '1') THEN
				OUTPUTSIGNAL <= OUTPUTSIGNAL + INPUT;
			END IF;
		END IF;
	END PROCESS;
		OUTPUT <= OUTPUTSIGNAL;
	
END DATAFLOW;