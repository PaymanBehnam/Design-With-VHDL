
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use work.my_pack.all;
entity routing is
end routing;

--}} End of automatically maintained section

architecture routing of routing is

begin
end routing;
